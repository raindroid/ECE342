module de1soc_top 
(
	// These are the board inputs/outputs required for all the ECE342 labs.
	// Each lab can use the subset it needs -- unused pins will be ignored.
	
    // Clock pins
    input                     CLOCK_50,

    // Seven Segment Displays
    output      [6:0]         HEX0,
    output      [6:0]         HEX1,
    output      [6:0]         HEX2,
    output      [6:0]         HEX3,
    output      [6:0]         HEX4,
    output      [6:0]         HEX5,

    // Pushbuttons
    input       [3:0]         KEY,

    // LEDs
    output      [9:0]         LEDR,

    // Slider Switches
    input       [9:0]         SW,

    // VGA
    output      [7:0]         VGA_B,
    output                    VGA_BLANK_N,
    output                    VGA_CLK,
    output      [7:0]         VGA_G,
    output                    VGA_HS,
    output      [7:0]         VGA_R,
    output                    VGA_SYNC_N,
    output                    VGA_VS
);

// This generates a one-time ACTIVE-LOW asynchronous reset
// signal on powerup. You can use it for the Qsys system.
logic reset_n;
logic [1:0] reset_reg;
always_ff @ (posedge CLOCK_50) begin
	reset_n <= reset_reg[0];
	reset_reg <= {1'b1, reset_reg[1]};
end

//
// INSTANTIATE QSYS SYSTEM HERE
//

// Implements a simple Nios II system for the DE-series board.
// Inputs:SW7−0 are parallel port inputs to the Nios II system CLOCK_50 is the system clock
//        KEY0 is the active-low system reset
//         LEDR7−0 are parallel port outputs from the Nios II system
// Outputs:
endmodule

module lights (CLOCK_50, SW, KEY, LEDR);
	input CLOCK_50; 
	input [7:0] SW; 
	input [0:0] KEY; 
	output [7:0] LEDR;
// Instantiate the Nios II system module generated by the Qsys tool: 
	nios_system NiosII (.clk_clk(CLOCK_50), 
							  .reset_reset_n(KEY), 
							  .switches_export(SW), 
							  .leds_export(LEDR));
endmodule


