//REVIEW  CPU moduls

module cpu (
    input clk,
    input reset,

    output logic [15:0] o_mem_addr,
    output logic        o_mem_rd,
    input[15:0]         o_mem_rddata,
    output logic        o_mem_wr,
    output logic [15:0] o_mem_wrdata
);

    // Datapath


    // Control FSM
    
endmodule