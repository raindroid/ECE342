/**
 * REVIEW 
 * module fast_adder
 */

module fast_adder_back #
(
    parameter N = 11    
)
(
    input [N-1:0] A,
    input [N-1:0] B,
    input Cin,

    output logic Cout,
    output logic [N - 1: 0]S
);

    logic [N-1: 0] g, p;
    logic [N: 0] C;

    genvar i;

    assign C[0] = Cin;
    assign Cout = C[N];

    // NOTE Connect g_i, p_i
    generate 
        for (i = 0; i < N; i++) begin : adder_units
            assign g[i] = A[i] & B[i];
            assign p[i] = A[i] | B[i];
            assign C[i + 1] = g[i] | (p[i] & C[i]);   // NOTE this is not exactly the same as CLA during the lecture
            assign S[i] =  A[i] ^ B[i] ^ C[i];
        end
    endgenerate


//     // REVIEW generated by WTM.py
//     logic [10: 0] ai, bi, gi, pi, si;
//     logic [11: 0] ci;

//     assign ai = A[10:0];
//     assign bi = B[10:0];
//     assign S = si[10:0];
//     assign ci[0] = Cin;
//     assign Cout = ci[N];

//     // NOTE connect all gi, pi, si
//     assign gi[0]        = ai[0] & bi[0];
//     assign pi[0]        = ai[0] | bi[0];
//     assign si[0]        = ai[0] ^ bi[0] ^ ci[0];
//     assign gi[1]        = ai[1] & bi[1];
//     assign pi[1]        = ai[1] | bi[1];
//     assign si[1]        = ai[1] ^ bi[1] ^ ci[1];
//     assign gi[2]        = ai[2] & bi[2];
//     assign pi[2]        = ai[2] | bi[2];
//     assign si[2]        = ai[2] ^ bi[2] ^ ci[2];
//     assign gi[3]        = ai[3] & bi[3];
//     assign pi[3]        = ai[3] | bi[3];
//     assign si[3]        = ai[3] ^ bi[3] ^ ci[3];
//     assign gi[4]        = ai[4] & bi[4];
//     assign pi[4]        = ai[4] | bi[4];
//     assign si[4]        = ai[4] ^ bi[4] ^ ci[4];
//     assign gi[5]        = ai[5] & bi[5];
//     assign pi[5]        = ai[5] | bi[5];
//     assign si[5]        = ai[5] ^ bi[5] ^ ci[5];
//     assign gi[6]        = ai[6] & bi[6];
//     assign pi[6]        = ai[6] | bi[6];
//     assign si[6]        = ai[6] ^ bi[6] ^ ci[6];
//     assign gi[7]        = ai[7] & bi[7];
//     assign pi[7]        = ai[7] | bi[7];
//     assign si[7]        = ai[7] ^ bi[7] ^ ci[7];
//     assign gi[8]        = ai[8] & bi[8];
//     assign pi[8]        = ai[8] | bi[8];
//     assign si[8]        = ai[8] ^ bi[8] ^ ci[8];
//     assign gi[9]        = ai[9] & bi[9];
//     assign pi[9]        = ai[9] | bi[9];
//     assign si[9]        = ai[9] ^ bi[9] ^ ci[9];
//     assign gi[10]       = ai[10] & bi[10];
//     assign pi[10]       = ai[10] | bi[10];
//     assign si[10]       = ai[10] ^ bi[10] ^ ci[10];

//     // NOTE connect all ci
//     assign ci[1] = ci[0] & pi[0] | gi[0];
//     assign ci[2] = ci[0] & pi[0] & pi[1] | gi[0] & pi[1] | gi[1];
//     assign ci[3] = ci[0] & pi[0] & pi[1] & pi[2] | gi[0] & pi[1] & pi[2] | gi[1] & pi[2] | gi[2];
//     assign ci[4] = ci[0] & pi[0] & pi[1] & pi[2] & pi[3] | gi[0] & pi[1] & pi[2] & pi[3] | gi[1] & pi[2] & pi[3] | gi[2] & pi[3] | gi[3];
//     assign ci[5] = ci[0] & pi[0] & pi[1] & pi[2] & pi[3] & pi[4] | gi[0] & pi[1] & pi[2] & pi[3] & pi[4] | gi[1] & pi[2] & pi[3] & pi[4] | gi[2] & pi[3] & pi[4] | gi[3] & pi[4] | gi[4];
//     assign ci[6] = ci[0] & pi[0] & pi[1] & pi[2] & pi[3] & pi[4] & pi[5] | gi[0] & pi[1] & pi[2] & pi[3] & pi[4] & pi[5] | gi[1] & pi[2] & pi[3] & pi[4] & pi[5] | gi[2] & pi[3] & pi[4] & pi[5] | gi[3] & pi[4] & pi[5] | gi[4] & pi[5] | gi[5];
//     assign ci[7] = ci[0] & pi[0] & pi[1] & pi[2] & pi[3] & pi[4] & pi[5] & pi[6] | gi[0] & pi[1] & pi[2] & pi[3] & pi[4] & pi[5] & pi[6] | gi[1] & pi[2] & pi[3] & pi[4] & pi[5] & pi[6] | gi[2] & pi[3] & pi[4] & pi[5] & pi[6] | gi[3] & pi[4] & pi[5] & pi[6] | gi[4] & pi[5] & pi[6] | gi[5] & pi[6] | gi[6];
//     assign ci[8] = ci[0] & pi[0] & pi[1] & pi[2] & pi[3] & pi[4] & pi[5] & pi[6] & pi[7] | gi[0] & pi[1] & pi[2] & pi[3] & pi[4] & pi[5] & pi[6] & pi[7] | gi[1] & pi[2] & pi[3] & pi[4] & pi[5] & pi[6] & pi[7] | gi[2] & pi[3] & pi[4] & pi[5] & pi[6] & pi[7] | gi[3] & pi[4] & pi[5] & pi[6] & pi[7] | gi[4] & pi[5] & pi[6] & pi[7] | gi[5] & pi[6] & pi[7] | gi[6] & pi[7] | gi[7];
//     assign ci[9] = ci[0] & pi[0] & pi[1] & pi[2] & pi[3] & pi[4] & pi[5] & pi[6] & pi[7] & pi[8] | gi[0] & pi[1] & pi[2] & pi[3] & pi[4] & pi[5] & pi[6] & pi[7] & pi[8] | gi[1] & pi[2] & pi[3] & pi[4] & pi[5] & pi[6] & pi[7] & pi[8] | gi[2] & pi[3] & pi[4] & pi[5] & pi[6] & pi[7] & pi[8] | gi[3] & pi[4] & pi[5] & pi[6] & pi[7] & pi[8] | gi[4] & pi[5] & pi[6] & pi[7] & pi[8] | gi[5] & pi[6] & pi[7] & pi[8] | gi[6] & pi[7] & pi[8] | gi[7] & pi[8] | gi[8];
//     assign ci[10] = ci[0] & pi[0] & pi[1] & pi[2] & pi[3] & pi[4] & pi[5] & pi[6] & pi[7] & pi[8] & pi[9] | gi[0] & pi[1] & pi[2] & pi[3] & pi[4] & pi[5] & pi[6] & pi[7] & pi[8] & pi[9] | gi[1] & pi[2] & pi[3] & pi[4] & pi[5] & pi[6] & pi[7] & pi[8] & pi[9] | gi[2] & pi[3] & pi[4] & pi[5] & pi[6] & pi[7] & pi[8] & pi[9] | gi[3] & pi[4] & pi[5] & pi[6] & pi[7] & pi[8] & pi[9] | gi[4] & pi[5] & pi[6] & pi[7] & pi[8] & pi[9] | gi[5] & pi[6] & pi[7] & pi[8] & pi[9] | gi[6] & pi[7] & pi[8] & pi[9] | gi[7] & pi[8] & pi[9] | gi[8] & pi[9] | gi[9];
//     assign ci[11] = ci[0] & pi[0] & pi[1] & pi[2] & pi[3] & pi[4] & pi[5] & pi[6] & pi[7] & pi[8] & pi[9] & pi[10] | gi[0] & pi[1] & pi[2] & pi[3] & pi[4] & pi[5] & pi[6] & pi[7] & pi[8] & pi[9] & pi[10] | gi[1] & pi[2] & pi[3] & pi[4] & pi[5] & pi[6] & pi[7] & pi[8] & pi[9] & pi[10] 
// | gi[2] & pi[3] & pi[4] & pi[5] & pi[6] & pi[7] & pi[8] & pi[9] & pi[10] | gi[3] & pi[4] & pi[5] & pi[6] & pi[7] & pi[8] & pi[9] & pi[10] | gi[4] & pi[5] & pi[6] & pi[7] & pi[8] & pi[9] & pi[10] | gi[5] & pi[6] & pi[7] & pi[8] & pi[9] & pi[10] | gi[6] & pi[7] & pi[8] & pi[9] & pi[10] 
// | gi[7] & pi[8] & pi[9] & pi[10] | gi[8] & pi[9] & pi[10] | gi[9] & pi[10] | gi[10];



endmodule