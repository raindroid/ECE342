// REVIEW line_drawing_algo module

    module line_drawing_algo (
        input clk,
        input reset,

        input i_start,
        input [8:0] i_x0,
        input [7:0] i_y0,
        input [8:0] i_x1,
        input [7:0] i_y1,
        input [2:0] i_color,

        output o_done,
        output 
    );
        
    endmodule